`timescale 1ns/1ps
module axi_lite_aphs
#(parameter
    C_S_AXI_ADDR_WIDTH = 8,    //the determinte the size of registers
    C_S_AXI_DATA_WIDTH = 32
)(
    input  wire                          ACLK,
    input  wire                          ARESET,
    input  wire                          ACLK_EN,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0] AWADDR,
    input  wire                          AWVALID,
    output wire                          AWREADY,
    input  wire [C_S_AXI_DATA_WIDTH-1:0] WDATA,
    input  wire [C_S_AXI_DATA_WIDTH/8-1:0] WSTRB,
    input  wire                          WVALID,
    output wire                          WREADY,
    output wire [1:0]                    BRESP,
    output wire                          BVALID,
    input  wire                          BREADY,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0] ARADDR,
    input  wire                          ARVALID,
    output wire                          ARREADY,
    output wire [C_S_AXI_DATA_WIDTH-1:0] RDATA,
    output wire [1:0]                    RRESP,
    output wire                          RVALID,
    input  wire                          RREADY,
    
    //ap_ctrl_hs bus
    output wire                          ap_start,
    input  wire                          ap_done,
    input  wire                          ap_ready,
    input  wire                          ap_idle,
    input  wire [0:0]                    ap_local_deadlock,
    output wire                          interrupt,
    
//   
    output wire [31:0]                   reg15_o,
    input  wire [31:0]                   reg15_i,
      
      output wire [31:0]                   reg14_o,
      input  wire [31:0]                   reg14_i,
      
      output wire [31:0]                   reg13_o,
      input  wire [31:0]                   reg13_i,
      
      output wire [31:0]                   reg12_o,
      input  wire [31:0]                   reg12_i,
      
      output wire [31:0]                   reg11_o,
      input  wire [31:0]                   reg11_i,
      
      output wire [31:0]                   reg10_o,
      input  wire [31:0]                   reg10_i,
      
      output wire [31:0]                   reg9_o,
      input  wire [31:0]                   reg9_i,
      
      output wire [31:0]                   reg8_o,
      input  wire [31:0]                   reg8_i,
      
      output wire [31:0]                   reg7_o,
      input  wire [31:0]                   reg7_i,
      
      output wire [31:0]                   reg6_o,
      input  wire [31:0]                   reg6_i,
      
      output wire [31:0]                   reg5_o,
      input  wire [31:0]                   reg5_i,
      
      output wire [31:0]                   reg4_o,
      input  wire [31:0]                   reg4_i,
      
      output wire [31:0]                   reg3_o,
      input  wire [31:0]                   reg3_i,
      
      output wire [31:0]                   reg2_o,
      input  wire [31:0]                   reg2_i,
      
      output wire [31:0]                   reg1_o,
      input  wire [31:0]                   reg1_i,
      
      output wire [31:0]                   reg0_o,
      input  wire [31:0]                   reg0_i
     
);
//------------------------Address Info-------------------
// 0x00 : Control signals
//        bit 0  - ap_start (Read/Write/COH)
//        bit 1  - ap_done (Read/COR)
//        bit 2  - ap_idle (Read)
//        bit 3  - ap_ready (Read/COR)
//        bit 7  - auto_restart (Read/Write)
//        others - reserved
// 0x04 : Global Interrupt Enable Register
//        bit 0  - Global Interrupt Enable (Read/Write)
//        others - reserved
// 0x08 : IP Interrupt Enable Register (Read/Write)
//        bit 0 - enable ap_done interrupt (Read/Write)
//        bit 1 - enable ap_ready interrupt (Read/Write)
//        bit 5 - enable ap_local_deadlock interrupt (Read/Write)
//        others - reserved
// 0x0c : IP Interrupt Status Register (Read/TOW)
//        bit 0 - ap_done (COR/TOW)
//        bit 1 - ap_ready (COR/TOW)
//        bit 5 - ap_local_deadlock (COR/TOW)
//        others - reserved

// (SC = Self Clear, COR = Clear on Read, TOW = Toggle on Write, COH = Clear on Handshake)

//------------------------Parameter----------------------
localparam
    ADDR_AP_CTRL           = 8'h00,
    ADDR_GIE               = 8'h04,
    ADDR_IER               = 8'h08,
    ADDR_ISR               = 8'h0c,
    //the bk lite interface
     ADDR_REG15             = 8'h4C,
     ADDR_REG14             = 8'h48,
     ADDR_REG13             = 8'h44,
     ADDR_REG12             = 8'h40,
     ADDR_REG11             = 8'h3C,
     ADDR_REG10             = 8'h38,
     ADDR_REG9              = 8'h34,
     ADDR_REG8              = 8'h30,
     ADDR_REG7              = 8'h2c,
     ADDR_REG6              = 8'h28,
     ADDR_REG5              = 8'h24,
     ADDR_REG4              = 8'h20,
     ADDR_REG3              = 8'h1C,
     ADDR_REG2              = 8'h18,
    ADDR_REG1              = 8'h14,
    ADDR_REG0              = 8'h10,
    
    
    
    WRIDLE                 = 2'd0,
    WRDATA                 = 2'd1,
    WRRESP                 = 2'd2,
    WRRESET                = 2'd3,
    RDIDLE                 = 2'd0,
    RDDATA                 = 2'd1,
    RDRESET                = 2'd2,
    ADDR_BITS                = 9;   //512 address

//------------------------Local signal-------------------
    reg  [1:0]                    wstate = WRRESET;
    reg  [1:0]                    wnext;
    reg  [ADDR_BITS-1:0]          waddr;
    wire [C_S_AXI_DATA_WIDTH-1:0] wmask;
    wire                          aw_hs;
    wire                          w_hs;
    reg  [1:0]                    rstate = RDRESET;
    reg  [1:0]                    rnext;
    reg  [C_S_AXI_DATA_WIDTH-1:0] rdata;
    wire                          ar_hs;
    wire [ADDR_BITS-1:0]          raddr;
    // internal registers
    reg                           int_ap_idle;
    reg                           int_ap_ready = 1'b0;
    wire                          task_ap_ready;
    reg                           int_ap_done = 1'b0;
    wire                          task_ap_done;
    reg                           int_task_ap_done = 1'b0;
    reg                           int_ap_start = 1'b0;
    reg                           int_auto_restart = 1'b0;
    reg                           auto_restart_status = 1'b0;
    wire                          auto_restart_done;
    reg                           int_gie = 1'b0;
    reg  [5:0]                    int_ier = 6'b0;
    reg  [5:0]                    int_isr = 6'b0;
    
//the bk lite interface    
    reg  [31:0]                   int_reg15 = 'b0;
    reg  [31:0]                   int_reg14 = 'b0;
    reg  [31:0]                   int_reg13 = 'b0;
    reg  [31:0]                   int_reg12 = 'b0;
    reg  [31:0]                   int_reg11 = 'b0;
    reg  [31:0]                   int_reg10 = 'b0;
    reg  [31:0]                   int_reg9 = 'b0;
    reg  [31:0]                   int_reg8 = 'b0;
    reg  [31:0]                   int_reg7 = 'b0;
    reg  [31:0]                   int_reg6 = 'b0;
    reg  [31:0]                   int_reg5 = 'b0;
    reg  [31:0]                   int_reg4 = 'b0;
    reg  [31:0]                   int_reg3 = 'b0;
    reg  [31:0]                   int_reg2 = 'b0;
    reg  [31:0]                   int_reg1 = 'b0;
    reg  [31:0]                   int_reg0 = 'b0;

//------------------------Instantiation------------------


//------------------------AXI write fsm------------------
assign AWREADY = (wstate == WRIDLE);
assign WREADY  = (wstate == WRDATA);
assign BRESP   = 2'b00;  // OKAY
assign BVALID  = (wstate == WRRESP);
assign wmask   = { {8{WSTRB[3]}}, {8{WSTRB[2]}}, {8{WSTRB[1]}}, {8{WSTRB[0]}} };
assign aw_hs   = AWVALID & AWREADY;
assign w_hs    = WVALID & WREADY;

// wstate
always @(posedge ACLK) begin
    if (ARESET)
        wstate <= WRRESET;
    else if (ACLK_EN)
        wstate <= wnext;
end

// wnext
always @(*) begin
    case (wstate)
        WRIDLE:
            if (AWVALID)
                wnext = WRDATA;
            else
                wnext = WRIDLE;
        WRDATA:
            if (WVALID)
                wnext = WRRESP;
            else
                wnext = WRDATA;
        WRRESP:
            if (BREADY)
                wnext = WRIDLE;
            else
                wnext = WRRESP;
        default:
            wnext = WRIDLE;
    endcase
end

// waddr
always @(posedge ACLK) begin
    if (ACLK_EN) begin
        if (aw_hs)
            waddr <= AWADDR[ADDR_BITS-1:0];
    end
end

//------------------------AXI read fsm-------------------
assign ARREADY = (rstate == RDIDLE);
assign RDATA   = rdata;
assign RRESP   = 2'b00;  // OKAY
assign RVALID  = (rstate == RDDATA);
assign ar_hs   = ARVALID & ARREADY;
assign raddr   = ARADDR[ADDR_BITS-1:0];

// rstate
always @(posedge ACLK) begin
    if (ARESET)
        rstate <= RDRESET;
    else if (ACLK_EN)
        rstate <= rnext;
end

// rnext
always @(*) begin
    case (rstate)
        RDIDLE:
            if (ARVALID)
                rnext = RDDATA;
            else
                rnext = RDIDLE;
        RDDATA:
            if (RREADY & RVALID)
                rnext = RDIDLE;
            else
                rnext = RDDATA;
        default:
            rnext = RDIDLE;
    endcase
end

// rdata
always @(posedge ACLK) begin
    if (ACLK_EN) begin
        if (ar_hs) begin
            rdata <= 'b0;
            case (raddr)
                ADDR_AP_CTRL: begin
                    rdata[0] <= int_ap_start;
                    rdata[1] <= int_task_ap_done;
                    rdata[2] <= int_ap_idle;
                    rdata[3] <= int_ap_ready;
                    rdata[7] <= int_auto_restart;
                end
                ADDR_GIE: begin
                    rdata <= int_gie;
                end
                ADDR_IER: begin
                    rdata <= int_ier;
                end
                ADDR_ISR: begin
                    rdata <= int_isr;
                end

                 ADDR_REG15: begin
                     rdata <= int_reg15;
                 end
                 ADDR_REG14: begin
                     rdata <= int_reg14;
                 end
                 ADDR_REG13: begin
                     rdata <= int_reg13;
                 end
                 ADDR_REG12: begin
                     rdata <= int_reg12;
                 end
                 ADDR_REG11: begin
                     rdata <= int_reg11;
                 end
                 ADDR_REG10: begin
                     rdata <= int_reg10;
                 end
                 ADDR_REG9: begin
                     rdata <= int_reg9;
                 end
                 ADDR_REG8: begin
                     rdata <= int_reg8;
                 end
                 ADDR_REG7: begin
                     rdata <= int_reg7;
                 end
                 ADDR_REG6: begin
                     rdata <= int_reg6;
                 end
                 ADDR_REG5: begin
                     rdata <= int_reg5;
                 end
                 ADDR_REG4: begin
                     rdata <= int_reg4;
                 end
                 ADDR_REG3: begin
                     rdata <= int_reg3;
                 end
                 ADDR_REG2: begin
                     rdata <= int_reg2;
                 end
                ADDR_REG1: begin
                    rdata <= int_reg1;
                end
                ADDR_REG0: begin
                    rdata <= int_reg0;
                end
               
            endcase
        end
    end
end


//------------------------Register logic-----------------
assign interrupt         = int_gie & (|int_isr);
assign ap_start          = int_ap_start;
assign task_ap_done      = (ap_done && !auto_restart_status) || auto_restart_done;
assign task_ap_ready     = ap_ready && !int_auto_restart;
assign auto_restart_done = auto_restart_status && (ap_idle && !int_ap_idle);

         assign reg15_o   = int_reg15;
         assign reg14_o   = int_reg14;
         assign reg13_o   = int_reg13;
         assign reg12_o   = int_reg12;
         assign reg11_o   = int_reg11;
         assign reg10_o   =  int_reg10;
         assign reg9_o    = int_reg9;
         assign reg8_o    = int_reg8;
         assign reg7_o    = int_reg7;
         assign reg6_o    = int_reg6;
         assign reg5_o    = int_reg5;
         assign reg4_o    = int_reg4;
         assign reg3_o    = int_reg3;
         assign reg2_o    = int_reg2;
         assign reg1_o    = int_reg1;
         assign reg0_o    = int_reg0;


// int_ap_start
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_start <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_AP_CTRL && WSTRB[0] && WDATA[0])
            int_ap_start <= 1'b1;
        else if (ap_ready)
            int_ap_start <= int_auto_restart; // clear on handshake/auto restart
    end
end

// int_ap_done
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_done <= 1'b0;
    else if (ACLK_EN) begin
            int_ap_done <= ap_done;
    end
end

// int_task_ap_done
always @(posedge ACLK) begin
    if (ARESET)
        int_task_ap_done <= 1'b0;
    else if (ACLK_EN) begin
        if (task_ap_done)
            int_task_ap_done <= 1'b1;
        else if (ar_hs && raddr == ADDR_AP_CTRL)
            int_task_ap_done <= 1'b0; // clear on read
    end
end

// int_ap_idle
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_idle <= 1'b0;
    else if (ACLK_EN) begin
            int_ap_idle <= ap_idle;
    end
end

// int_ap_ready
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_ready <= 1'b0;
    else if (ACLK_EN) begin
        if (task_ap_ready)
            int_ap_ready <= 1'b1;
        else if (ar_hs && raddr == ADDR_AP_CTRL)
            int_ap_ready <= 1'b0;
    end
end

// int_auto_restart
always @(posedge ACLK) begin
    if (ARESET)
        int_auto_restart <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_AP_CTRL && WSTRB[0])
            int_auto_restart <=  WDATA[7];
    end
end

// auto_restart_status
always @(posedge ACLK) begin
    if (ARESET)
        auto_restart_status <= 1'b0;
    else if (ACLK_EN) begin
        if (int_auto_restart)
            auto_restart_status <= 1'b1;
        else if (ap_idle)
            auto_restart_status <= 1'b0;
    end
end

// int_gie
always @(posedge ACLK) begin
    if (ARESET)
        int_gie <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_GIE && WSTRB[0])
            int_gie <= WDATA[0];
    end
end

// int_ier
always @(posedge ACLK) begin
    if (ARESET)
        int_ier <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_IER && WSTRB[0])
            int_ier <= WDATA[5:0];
    end
end

// int_isr[0]
always @(posedge ACLK) begin
    if (ARESET)
        int_isr[0] <= 1'b0;
    else if (ACLK_EN) begin
        if (int_ier[0] & ap_done)
            int_isr[0] <= 1'b1;
        else if (w_hs && waddr == ADDR_ISR && WSTRB[0])
            int_isr[0] <= int_isr[0] ^ WDATA[0]; // toggle on write
    end
end

// int_isr[1]
always @(posedge ACLK) begin
    if (ARESET)
        int_isr[1] <= 1'b0;
    else if (ACLK_EN) begin
        if (int_ier[1] & ap_ready)
            int_isr[1] <= 1'b1;
        else if (w_hs && waddr == ADDR_ISR && WSTRB[0])
            int_isr[1] <= int_isr[1] ^ WDATA[1]; // toggle on write
    end
end

// int_isr[5]
always @(posedge ACLK) begin
    if (ARESET)
        int_isr[5] <= 1'b0;
    else if (ACLK_EN) begin
        if (int_ier[5] & ap_local_deadlock)
            int_isr[5] <= 1'b1;
        else if (w_hs && waddr == ADDR_ISR && WSTRB[0])
            int_isr[5] <= int_isr[5] ^ WDATA[5]; // toggle on write
    end
end

/******************************************bk lite***************************************************************/
// int_reg15[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg15[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG15)
            int_reg15[31:0] <= (WDATA[31:0] & wmask) | reg15_i;
    end
end

// int_reg14[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg14[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG14)
            int_reg14[31:0] <= (WDATA[31:0] & wmask) |  reg14_i;
    end
end

// int_reg13[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg13[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG13)
            int_reg13[31:0] <= (WDATA[31:0] & wmask) |  reg13_i ;
    end
end

// int_reg12[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg12[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG12)
            int_reg12[31:0] <= (WDATA[31:0] & wmask) |  reg12_i ;
    end
end
// int_reg11[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg11[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG11)
            int_reg11[31:0] <= (WDATA[31:0] & wmask) |  reg11_i ;
    end
end

// int_reg10[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg10[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG10)
            int_reg10[31:0] <= (WDATA[31:0] & wmask) | reg10_i ;
    end
end

// int_reg9[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg9[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG9)
            int_reg9[31:0] <= (WDATA[31:0] & wmask) | reg9_i ;
    end
end

// int_reg8[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg8[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG8)
            int_reg8[31:0] <= (WDATA[31:0] & wmask) | reg8_i ;
    end
end

// int_reg7[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg7[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG7)
            int_reg7[31:0] <= (WDATA[31:0] & wmask) | reg7_i ;
    end
end

// int_reg6[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg6[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG6)
            int_reg6[31:0] <= (WDATA[31:0] & wmask) | reg6_i ;
    end
end

// int_reg5[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg5[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG5)
            int_reg5[31:0] <= (WDATA[31:0] & wmask) | reg5_i ;
    end
end

// int_reg4[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg4[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG4)
            int_reg4[31:0] <= (WDATA[31:0] & wmask) | reg4_i ;
    end
end

// int_reg3[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg3[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG3)
            int_reg3[31:0] <= (WDATA[31:0] & wmask) | reg3_i ;
    end
end

// int_reg2[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg2[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG2)
            int_reg2[31:0] <= (WDATA[31:0] & wmask) | reg2_i ;
    end
end

// int_reg1[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg1[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG1)
            int_reg1[31:0] <= (WDATA[31:0] & wmask) | reg1_i ;
    end
end

// int_reg0[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_reg0[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_REG0)
            int_reg0[31:0] <= (WDATA[31:0] & wmask) | reg0_i ;
    end
end

//------------------------Memory logic-------------------

endmodule